��S w e d i s h  
 [ 1 1 1 ]  
 1 1 6 4 = B e h a n d l a   h e l a   b i l d e n  
 1 1 6 2 = N o l l s t � l l  
 1 1 6 3 = H j � l p  
 [ 1 1 5 ]  
 0 = C o d e c s  
 1 2 8 3 = C o d e c s   s o m   s t � d s  
 1 0 1 1 = X V I D  
 1 0 1 7 = A n v � n d   X v i D  
 1 0 1 2 = D i v X   3  
 1 0 1 3 = D i v X   4  
 1 0 1 6 = A n v � n d   X v i D  
 1 0 1 4 = D i v X   5  
 1 0 1 8 = A n v � n d   X v i D  
 1 0 5 0 = B L Z 0  
 1 0 1 9 = A n v � n d   X v i D  
 1 0 2 4 = M P 4 3  
 1 0 2 3 = M P 4 2  
 1 0 2 5 = M P 4 1  
 1 0 2 6 = W M V 1  
 1 0 4 8 = H . 2 6 3 +  
 1 0 4 9 = M P E G 1  
 1 0 5 3 = A n v � n d   L i b m p e g 2  
 1 0 5 2 = M P E G 2  
 1 0 5 4 = A n v � n d   L i b m p e g 2  
 1 0 5 5 = M J P E G  
 1 0 5 6 = D V  
 1 0 1 5 = R �   v i d e o  
 1 2 8 4 = F � r g r y m d e r   f � r   o u t p u t   s o m   s t � d s  
 1 0 2 0 = Y V 1 2  
 1 0 2 1 = Y U Y 2  
 1 0 2 2 = Y V Y U  
 1 0 2 7 = U Y V Y  
 1 0 5 1 = R G B 3 2  
 1 0 2 8 = R G B 2 4  
 1 0 2 9 = R G B 1 6  
 1 0 3 0 = R G B 1 5  
 1 0 3 1 = A n v � n d   o v e r l a y   m i x e r  
 1 1 6 6 = R e g i s t r e r a   i n t e   o m a r k e r a d e   c o d e c s  
 [ 1 1 6 ]  
 0 = I n f o r m a t i o n  
 1 2 8 4 = I n f o r m a t i o n  
 1 0 5 0 = N u   s p e l a s  
 1 0 5 5 = C o d e c  
 1 2 6 4 = F � r g r y m d   f � r   o u t p u t :  
 1 0 5 4 = D i m e n s i o n e r :  
 1 2 6 5 = F P S :  
 1 0 5 9 = N u v a r a n d e   r u t a :  
 1 2 6 6 = F P S   f � r   a v k o d a r e :  
 1 0 6 0 = B i t r a t e :  
 [ 1 3 2 ]  
 0 = T y p s n i t t  
 1 2 5 9 = T y p s n i t t  
 1 1 1 0 = S t o r l e k  
 1 1 1 6 = M e l l a n r u m  
 1 1 1 4 = T e c k e n  
 1 1 0 8 = S t y r k a  
 1 1 2 4 = F � r g  
 1 1 1 8 = S k u g g s t y r k a  
 1 1 3 0 = S k u g g s t o r l e k  
 [ 1 4 1 ]  
 0 = O S D  
 1 1 8 2 = O S D  
 1 1 1 0 = S t o r l e k  
 1 1 1 6 = M e l l a n r u m  
 1 1 1 4 = T e c k e n  
 1 1 0 8 = S t y r k a  
 1 1 2 4 = F � r g  
 1 1 1 8 = S k u g g s t y r k a  
 1 1 3 0 = S k u g g s t o r l e k  
 [ 1 3 6 ]  
 0 = T r a y   &   d i a l o g   i n s t � l l n i n g a r  
 1 2 5 7 = T r a y   i k o n  
 1 0 7 0 = V i s a   t r a y   i k o n  
 1 2 5 8 = K o n f i g u r a t i o n s d i a l o g  
 1 0 7 1 = � t e r s t � l l   p o s i t i o n  
 1 0 7 2 = V i s a   h j � l p t e x t e r  
 1 2 9 3 = S p r � k  
 [ 1 4 3 ]  
 0 = T a n g e n t b o r d s s t y r n i n g  
 1 2 0 2 = A k t i v e r a d  
 [ 1 1 9 ]  
 0 = B i l d i n s t � l l n i n g a r  
 1 2 7 8 = F � r i n s t � l l n i n g a r  
 1 0 1 6 = N y  
 1 1 5 6 = L � s   f r � n   f i l . . .  
 1 1 5 5 = S p a r a   t i l l   f i l . . .  
 1 0 4 5 = B y t   n a m n  
 1 0 4 4 = T a   b o r t  
 1 0 5 1 = A u t o m a t i s k   i n l a d d n i n g  
 1 0 8 0 = F � r s � k   l a d d a   f � r i n s t � l l n i n g   f r � n   f i l   f � r s t  
 1 1 5 7 = R e g l e r   f � r   a u t o m a t i s k   i n l a d d n i n g  
 [ 1 2 0 ]  
 0 = E f t e r b e h a n d l i n g  
 1 0 7 3 = E f t e r b e h a n d l i n g  
 1 0 2 7 = F � r i n s t � l l n i n g a r  
 1 0 0 8 = A u t o m a t i s k   k v a l i t e t s k o n t r o l l  
 1 0 2 8 = E g n a   i n s t � l l n i n g a r  
 1 2 7 0 = L u m i n a n s  
 1 2 7 1 = C h r o m a  
 1 2 7 2 = A v b l o c k n i n g   ( H )  
 1 2 7 3 = A v b l o c k n i n g   ( V )  
 1 2 7 4 = D e r i n g  
 1 1 5 8 = B e h a n d l i n g s s t y r k a  
 1 1 6 0 = B e h a n d l i n g s m e t o d :  
 1 2 3 8 = m p l a y e r  
 1 2 3 9 = N i c ' s  
 1 0 3 7 = T e m p o r a l t   b r u s f i l t e r  
 1 2 7 5 = N i v �   f i x  
 1 0 3 5 = L u m i n a n s  
 1 0 3 8 = H e l t   l u m a s p e c t r u m  
 1 0 3 6 = C h r o m a   ( e j   i m p l e m e n t e r a d )  
 1 2 4 2 = X   t r � s k e l  
 1 2 4 3 = Y   t r � s k e l  
 [ 1 2 5 ]  
 0 = B i l d e g e n s k a p e r  
 1 0 7 2 = B i l d e g e n s k a p e r  
 1 0 1 7 = L u m i n a n s � k n i n g  
 1 0 1 8 = L u m i n a n s o f f s e t  
 1 0 3 7 = G a m m a   k o r r i g e r i n g  
 1 0 2 5 = F � r g n y a n s  
 1 0 2 6 = F � r g m � t t n a d  
 [ 1 4 2 ]  
 0 = N i v � e r  
 1 1 7 0 = N i v � e r  
 1 1 7 9 = M o d i f i e r a   e n d a s t   l u m a  
 1 1 8 4 = V i s a   h i s t o g r a m  
 1 1 8 5 = H e l t   s p e c t r u m  
 1 2 9 1 = I n p u t  
 1 2 6 7 = O u t p u t  
 1 1 8 1 = G a m m a k o r r i g e r i n g  
 [ 1 2 6 ]  
 0 = B r u s  
 1 0 3 8 = B r u s  
 1 0 6 7 = G a m m a l   b r u s a l g o r i t m  
 1 0 6 8 = N y   b r u s a l g o r i t m   ( a v i h )  
 1 0 6 9 = m p l a y e r   b r u s  
 1 2 3 2 = G e n o m s n i t t  
 1 0 3 9 = U n i f o r m t   b r u s  
 1 2 3 1 = M � n s t e r  
 1 0 4 1 = S t y r k a   p �   l u m i n a n s b r u s  
 1 0 4 9 = S t y r k a   p �   c h r o m a b r u s  
 [ 1 2 7 ]  
 0 = S k � r p a  
 1 0 6 5 = S k � r p a  
 1 0 6 3 = x s k � r p a  
 1 0 6 4 = a v s k � r p n i n g s m a s k  
 1 0 6 6 = m s k � r p a  
 1 2 1 6 = h � g   k v a l i t e t  
 1 2 1 5 = b a r a   m a s k  
 1 0 6 7 = w a r p s k � r p a  
 1 0 1 9 = S t y r k a  
 1 0 2 1 = T r � s k e l  
 [ 1 2 8 ]  
 0 = B l u r   &   B R  
 1 1 3 4 = B l u r   & &   b r u s   r e d u c e r i n g  
 1 1 3 6 = S o f t e n  
 1 1 3 7 = T e m p o r a l u t j � m n i n g  
 1 2 3 2 = B e h a n d l a   f � r g  
 1 1 3 8 = L u m a u t j � m n a r e  
 1 1 3 9 = C h r o m i n a n c e u t j � m n a r e  
 1 1 4 0 = G r a d u a l   a v b r u s n i n g  
 [ 1 3 7 ]  
 0 = O f f s e t  
 1 1 4 8 = O f f s e t  
 1 1 4 9 = L u m a   o f f s e t   X  
 1 1 5 1 = L u m a   o f f s e t   Y  
 1 1 5 3 = C h r o m a   o f f s e t   X  
 1 1 2 0 = C h r o m a   o f f s e t   Y  
 [ 1 3 9 ]  
 0 = V i s a   R V  
 1 0 7 4 = V i s a   r � r e l s e v e k t o r e r  
 [ 1 7 2 ]  
 0 = F � n g a  
 1 2 1 6 = F � n g a  
 1 2 2 3 = V a r j e   r u t a  
 1 2 2 4 = E n   r u t a  
 1 2 2 6 = I n t e r v a l l  
 1 1 8 3 = P a t h  
 1 2 1 8 = . . .  
 1 2 6 1 = N a m n p r e f i x  
 1 2 6 3 = S i f f r o r   f � r   b i l d n u m r e r i n g  
 1 2 6 2 = B i l d f o r m a t  
 1 2 2 8 = F � n g a   n u  
 1 2 3 0 = K v a l i t e t  
 [ 1 1 3 ]  
 0 = T e x t n i n g  
 1 1 0 5 = T e x t n i n g  
 1 1 3 3 = S � k  
 1 1 8 3 = F i l  
 1 1 2 0 = . . .  
 1 1 2 2 = H o r i s o n t e l l   p o s i t i o n  
 1 1 2 6 = V e r t i k a l   p o s i t i o n  
 1 2 8 0 = F � r d r � j  
 1 2 8 1 = F a r t  
 1 2 4 4 = L a d d a   o m  
 1 1 2 4 = . . .  
 1 2 7 9 = S � k   i  
 [ 1 3 3 ]  
 0 = S t o r l e k   &   A s p e k t  
 1 0 8 3 = � n d r a   s t o r l e k  
 1 1 8 5 = S p e c i f i c e r a   s t o r l e k  
 1 2 8 5 = N y   s t o r l e k  
 1 1 8 6 = S p e c i f i c e r a   a s p e k t   r a t i o  
 1 2 8 6 = A s p e k t  
 1 1 8 7 = U t � k a   t i l l   n � s t a   m u l t i p e l   a v  
 1 1 8 9 = � n d r a   s t o r l e k   o m   . . .  
 1 2 8 7 = x  
 1 1 9 0 = o c h  
 1 2 8 8 = y  
 1 1 9 1 = � n d r a   s t o r l e k   o m   a n t a l e t   p u n k t e r  
 1 1 9 2 = s t � r r e   � n  
 1 1 8 8 = � n d r a   a l l t i d  
 1 2 8 9 = A s p e k t   r a t i o  
 1 1 0 0 = I n g e n   k o r r i g e r i n g   a v   a s p e k t   r a t i o  
 1 1 0 1 = B e h � l l   u r s p r u n g l i g   a s p e k t   r a t i o  
 1 1 0 2 = S � t t   a s p e k t   r a t i o   m a n u e l l t  
 1 2 9 0 = S v a r t a   k a n t e r  
 1 2 0 1 = H o r i s o n t e l l  
 1 2 0 0 = V e r t i k a l  
 1 1 9 9 = L � s  
 1 2 3 4 = O v e r l a y   a s p e k t   r a t i o :  
 [ 1 3 8 ]  
 0 = I n s t � l l n i n g a r  
 1 2 8 2 = S t o r l e k s i n s t � l l n i n g a r  
 1 2 8 5 = M e t o d  
 1 0 9 8 = L u m a   g a u s s i s k   b l u r  
 1 0 9 9 = C h r o m a   g a u s s i s k   b l u r  
 1 0 1 9 = L u m a s k � r p a  
 1 0 2 0 = C h r o m a s k � r p a  
 1 0 2 1 = P a r a m e t e r  
 [ 1 3 4 ]  
 0 = B e s k � r n i n g  
 1 1 3 7 = B e s k � r n i n g   & &   z o o m  
 1 1 3 8 = Z o o m  
 1 1 3 9 = B e s k � r n i n g  
 1 1 0 5 = H o r i s o n t e l l   f � r s t o r i n g  
 1 1 0 7 = V e r t i k a l   f � r s t o r i n g  
 1 1 4 0 = L � s  
 1 2 5 2 = T o p p  
 1 2 5 4 = V �  
 1 2 5 5 = H �  
 1 2 5 6 = B o t t e n  
 1 1 4 1 = P a n   & &   s c a n  
 1 1 0 9 = Z o o m  
 1 1 1 1 = H o r i s o n t e l l   p o s i t i o n  
 1 1 1 3 = V e r t i k a l   p o s i t i o n  
 [ 1 4 0 ]  
 0 = D e i n t e r l a c i n g  
 1 1 6 7 = D e i n t e r l a c i n g  
 1 1 6 9 = L i n j � r   i n t e r p o l e r i n g  
 1 1 7 0 = L i n j � r   b l a n d n i n g  
 1 1 7 1 = K u b i s k   i n t e r p o l e r i n g  
 1 1 7 3 = K u b i s k   b l a n d n i n g  
 1 1 7 2 = M e d i a n  
 1 1 7 4 = T o m s M o C o m p  
 1 2 0 7 = S � k s t y r k a :  
 1 2 0 9 = V � x l a   f � l t  
 1 1 7 5 = B o b   ( ? )  
 [ 1 7 3 ]  
 0 = O v e r l a y  
 1 2 3 5 = O v e r l a y k o n t r o l l  
 1 2 3 6 = L j u s s t y r k a  
 1 1 3 7 = K o n t r a s t  
 1 1 3 8 = F � r g n y a n s  
 1 1 3 9 = F � r g m � t t n a d  
 1 1 4 0 = S k � r p a  
 1 1 4 1 = G a m m a  
 [ 1 1 8 ]  
 0 = D i v e r s e  
 1 2 8 3 = D i v e r s e  
 1 0 1 6 = V � n d   b i l d  
 1 0 4 5 = I D C T  
 1 2 6 8 = V i d e o f � r d r � j n i n g :  
 1 2 6 9 = m s  
 1 0 4 7 = W o r k a r o u n d   e n c o d e r   b u g  
 1 2 9 4 = D e c i m e r i n g   a v   r a t i o  
 [ 1 0 2 ]  
 0 = O m  
 1 2 5 1 = f f d s h o w   M P E G - 4   V I D E O   A V K O D A R E  
 1 0 7 2 = D i r e c t S h o w   f i l t e r   b u i l d   d a t u m :  
 1 0 7 1 = l i b a v c o d e c   v e r s i o n  
 1 0 7 3 = x v i d   v e r s i o n  
  
  
  
  
 